`define BLACK       12'b0000_0000_0000
module vga(
        input clk,               // 100MHz
        input lcd_rst,             // 复位信号
        input select,            // 模式选择
        output hsync,            // 行同步信号
        output vsync,            // 场同步信号
        output [3:0] vga_r,      // VGA红色信号
        output [3:0] vga_g,      // VGA绿色信号
        output [3:0] vga_b       // VGA蓝色信号
    );

    // 行和列计数
    reg [9:0] x_cnt;
    reg [9:0] y_cnt;
    reg clk_vga = 0;
    reg clk_cnt = 0;

    // 生成25MHz VGA时钟
    always @(posedge clk) begin
        if (!lcd_rst)
            clk_vga <= 0;
        else if (clk_cnt == 1) begin
            clk_vga <= ~clk_vga;
            clk_cnt <= 0;
        end
        else
            clk_cnt <= clk_cnt + 1;
    end

    // VGA行和列计数
    always @ (posedge clk_vga) begin
        if (!lcd_rst)
            x_cnt <= 10'd0;
        else if (x_cnt == 10'd799)
            x_cnt <= 10'd0;
        else
            x_cnt <= x_cnt + 1;
    end

    always @ (posedge clk_vga) begin
        if (!lcd_rst)
            y_cnt <= 10'd0;
        else if (x_cnt == 10'd799) begin
            if (y_cnt == 10'd524)
                y_cnt <= 10'd0;
            else
                y_cnt <= y_cnt + 1;
        end
    end

    // VGA同步信号生成
    reg hsync_r, vsync_r;
    always @ (posedge clk_vga) begin
        if (!lcd_rst)
            hsync_r <= 1'b1;
        else if (x_cnt == 10'd0)
            hsync_r <= 1'b0;
        else if (x_cnt == 10'd96)
            hsync_r <= 1'b1;
    end

    always @ (posedge clk_vga) begin
        if (!lcd_rst)
            vsync_r <= 1'b1;
        else if (y_cnt == 10'd0)
            vsync_r <= 1'b0;
        else if (y_cnt == 10'd2)
            vsync_r <= 1'b1;
    end

    assign hsync = hsync_r;
    assign vsync = vsync_r;

    // 定义图案数据
    //XUPT logo  512X256
    parameter
        char_line0  = 512'h000000000000000000007FF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line1  = 512'h0000000000000000007FFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line2  = 512'h00000000000000000FFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line3  = 512'h00000000000000007FFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line4  = 512'h0000000000000003FFF800007FFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line5  = 512'h000000000000001FFE00000003FFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line6  = 512'h000000000000007FE0000000003FF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line7  = 512'h00000000000001FF000009800007FE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line8  = 512'h00000000000007FC0007FFC38000FF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line9  = 512'h0000000000001FE000EDF7C382003FC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line10 = 512'h0000000000003F800DB7B7CFE7C007F0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line11 = 512'h000000000000FE003F1CF7CDE37803FC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line12 = 512'h000000000001FC003797B987E33E00FE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line13 = 512'h000000000007F00718F00000067FC03F000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line14 = 512'h00000000000FC01B0C00000003D3101FC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line15 = 512'h00000000001F806F1801FFFE007F1C07E00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line16 = 512'h00000000003F00FE003FFFFFE00EB603F00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line17 = 512'h00000000007C018B01FFFFFFFE03FA01F80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line18 = 512'h0000000000F801880FFE0003FF80F3C0FC0000000000000000000000000000000000000000000000000000000000000000000000000000000000040000000000,
        char_line19 = 512'h0000000001F018F83FE000001FF03E607E00000000000000000000000000000000000000000000000000000000000000000000000000000000001E0000000000,
        char_line20 = 512'h0000000003E01800FF00000003FC04603F00000000000000000000000000000000000000000000000000000000000000000000000000000000003E0000000000,
        char_line21 = 512'h0000000007C07803F8000000007E073C1F8000000000000000000000000000000000000000003000000000000000C000000000000000000000003E0000000000,
        char_line22 = 512'h000000000F80FF07E0000000001F83E40FC00000000000000000000000000001E00000000000FC00000000000007FC00000000000000000000003E0000000000,
        char_line23 = 512'h000000001F81861F800000000007C0C607C00000000000000000000000000001F00000000003FF0000000000003FFE00000000000000000000303E0000000000,
        char_line24 = 512'h000000001F03E03E000000000003F0FD83E00000000000000000000000000001F8000000000FFF800000000000FFFE00000000070000000000F87E0000000000,
        char_line25 = 512'h000000003E07387C01FF0007FE00F83B81F000000000000001E0000000000003FC00000001FFFF80000000003FFFFC000000000F8000000000FCFC0700000000,
        char_line26 = 512'h000000007C0790F00FFFE03FFFC07C1F01F00000000000003FF8000000000003FE00000003FFFF00000000003FFFF0000000000FC000000000FFF81F00000000,
        char_line27 = 512'h000000007C0DE1E03FFFF87FFFF03E1FE0F8000000000003FFFC000000000C07FE00000000FFCF80000000001FFFCE000000000FE000000020FFF07F00000000,
        char_line28 = 512'h00000000F813C3C0FFFFFDFFFFF81F0FE07C0000000000FFFFFC000000001E07FC00000000FFFF80000000000FFFFFFFF800000FF000000070FFF1FE00000000,
        char_line29 = 512'h00000000F01C8781FFFFFFFFFFFC0F87107C0000000003FFFFFC000000001F0FFC00000001FFFF80007F8000007FFFFFFC00000FF00000007CFEFFFC00000000,
        char_line30 = 512'h00000001F0338F03FFFFFFFFFFFE07C2F03C0000000007FFFFF8000000001F8FF3C0000003FFFE0603FF800007FFFF9FFC00000FF00000003FFDFFF800000000,
        char_line31 = 512'h00000001F07B1F03FFFFFFFFFFFF03C3E03E000000000FFFFF80000000001F9FFFC000003FFFFF0F8FFE001E0FFFF83FFC00000FE00000003FFFFFF000000000,
        char_line32 = 512'h00000003E05E1E07FFFFFFFFFFFF81E0FC1E000000001FFFFF00000000001F9FFFC000003FFFFF1FFFFC003F1FFFFBFFF000001FC01C00003FFFFFE000000000,
        char_line33 = 512'h00000003E0FC3C0FFFFFFFFFFFFF80E0FC1F000000000FFFFFF0000000003F3FFFC000003FFFFF9FFFF8007FFFFFFBFFC000001FC1FF00003EFFFFE000000000,
        char_line34 = 512'h00000003C0CC3C0FFFFFFFFFFFFFC0F0E61F0000000003FFCFF0000000003F7F9FC000001FFF9FDFFFF0007FFFFE7C000000001FFFFF00003EFFFFC000000000,
        char_line35 = 512'h00000007C1EC780FFFFFFFFFFFFFC0703E0F0000000003FF0FF8000000003FFF3FC000000FEFFFBFFFE0007E1FFFFC000000001FFFFF00001EFFFFFFE0000000,
        char_line36 = 512'h00000007C1FC780FFFFFFFFFFFFFC078600F8000000003FF07FC1E0000007FFFFFC0000007FFFF7FDFC0007E1FFFE000000007FFFFFF00003EFFFFFFFC000000,
        char_line37 = 512'h0000000781F8F00FFFFFFFFFC3FFC0386F0F8000000001FF07FFFF800000FFFFFC00000007FFFE7FFF0000FE1F7C00000003FFFFFFFC0000FFFFFFFFFC000000,
        char_line38 = 512'h0000000F8398F00FFFE01FFF07FFC03C390F8000000001FF8FFFFFC00000FFFEE0000000FFFFF87FFE0000FC1EFC00000007FFFFFE000003EFFFE07FFC000000,
        char_line39 = 512'h0000000F80E0E00FFF800FFC1FFFC03C3F078000000001FFFFFC3FC00001FFFC0003C001FFFF7FBFFC0000FC7CFFFE00000FFFFFC000000FFFE7800000000000,
        char_line40 = 512'h0000000F83F1E00FFE0001F03FFF803C3707C000000001FFFFF87FC00001FDF87CFFE000FFEFFE3FFC000078E1FFFE00000FFFFFE000001FFF9E0F8000000000,
        char_line41 = 512'h0000000F83E1E007FFC00000FFFF801C1D07C000007C00FFFFF07FC0000063FFFFFFE00003EFFF3FFE000001E7FFFE000007F8FFF000001FFE7DFF8000000000,
        char_line42 = 512'h0000000F83F1E007FFFC0001FFFF001E3F87C00000FF01FFFFF0FFC000000FFFFFFFE00001DFFE3FFF000001EFFCFC00000301FBF800003FF0F7FF8000000000,
        char_line43 = 512'h0000000F03F1E003FFFF0003FFFE001E3F87C00000FF83FFFFE0FF800003FFFFFFFFC00001FFCE3FBF800003FC7CFC00000003F9FC00003FC3FFFF0000000000,
        char_line44 = 512'h0000000F03F1E001FFFFC003FFFC001E3E87C00000FFEFFFFFE1FE000FFFFFFFFE3FC00003FE1C3FCFC00003FFFFFC00000003F0FF00007F07F8FE0000000000,
        char_line45 = 512'h0000000F02E1C000FFFFE007FFF8001E1F07C00000FFFFFF9FC3F8001FFFFFFFFE078000FF8FFC3F8FC00003FFFFF800000007F07F80003C0FE3F80000000000,
        char_line46 = 512'h0000000F03B1C000FFFFF00FFFFC001E3187C000007FFFFF1FC3F0003FFFFF8FFE000007FC0FFC3F87E00003CFFCF80000000FE03FE000000F87FC0000000000,
        char_line47 = 512'h0000000F03F1E001FFFFF00FFFFE001E3187C000007FFFFF3F87E0003FFE3FFFF800003FF01FF83FC7E00001E7F9F00000000FC00FF800000F07FFFC00000000,
        char_line48 = 512'h0000000F03E1E003FFFFE00FFFFF001E3B87C000003FFFFF7F0FE0003FC01FFFC000003F803F003FF7F00001E3FFF00000003F8007FF00000007FFFE00000000,
        char_line49 = 512'h0000000F83F1E007FFFFC01FFFFF001E3C07C000001FFE7FFFFFC0000F000FFF0000001E01FC003FFFE00000E1FFE00000007F0003FFC00003FFFFFC00000000,
        char_line50 = 512'h0000000F8011E007FFFFC03FFFFF801C0F07C000000FFC3FFFFFC000000003FF8000000003F0003FFFE00000F7FFE0000000FE0000FFE0001FFFFE0000000000,
        char_line51 = 512'h0000000F83F0E00FFFFF80FFFFFF803C3F07C0000007FE7FFFFFC000000001FFE00000000FC0003F7FC00000FFFF8000000FFC00007FF0003FFFF80000000000,
        char_line52 = 512'h0000000F8300F00FFFFE03FFFFFFC03C220780000003FFFFFFFF8000000007FFFC000000FF80003F3FC000007FF0000000FFF800001FF8001FC1F80000000000,
        char_line53 = 512'h000000078000F00FFFFC0FFFFFFFC03C7B0F80000001FFFFFFFF800000001FE1FFE000007F00003F1F80000000F8000001FFF0000003F8000181F80000000000,
        char_line54 = 512'h00000007C138F00FFFFE7FFFFFFFC0787F0F80000000FFFFFFFF000000007F807FF000000C00003F02000000007E000001FFC000000070000003F80000000000,
        char_line55 = 512'h00000007C1F8780FFFFFFFFFFFFFC078460F80000000FFFFC0FC0000003FFF001FFC00000000003F00000000007FF30000FF0000000000000003F00000000000,
        char_line56 = 512'h00000007C16C780FFFFFFFFFFFFFC0F0FE0F000000007FFC01E00000007FFC0001FE00000000003E00000000003FFF8000F80000000000000007F00000000000,
        char_line57 = 512'h00000003E0FC3C0FFFFFFFFFFFFFC0F0FC1F000000003FE001800000007FE000003C00000000003E000000000007FF800000000000000000000FF00000000000,
        char_line58 = 512'h00000003E0CE3C07FFFFFFFFFFFF81E1F81F000000000FC000000000007F0000000000000000003E000000000000FF00000000000000000000FFE00000000000,
        char_line59 = 512'h00000003E0181E07FFFFFFFFFFFF81E1083E0000000000000000000000000000000000000000003E00000000000004000000000000000000FFFFC00000000000,
        char_line60 = 512'h00000001F03F0F03FFFFFFFFFFFF03C1D83E0000000000000000000000000000000000000000003E00000000000000000000000000000000FFFF800000000000,
        char_line61 = 512'h00000001F03F0F81FFFFFFFFFFFE0787F07C0000000000000000000000000000000000000000003C000000000000000000000000000000003FC0000000000000,
        char_line62 = 512'h00000000F808C7C0FFFFFFFFFFFC0F01C07C000000000000000000000000000000000000000000FC000000000000000000000000000000000000000000000000,
        char_line63 = 512'h00000000FC1FC3E07FFFFCFFFFF81F0FE0F8000000000000000000000000000000000000000000F8000000000000000000000000000000000000000000000000,
        char_line64 = 512'h000000007C0E61F03FFFF07FFFE03E1F00F800000000000000000000000000000000000000000030000000000000000000000000000000000000000000000000,
        char_line65 = 512'h000000003E07D0F80FFFC01FFF807C3DC1F000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line66 = 512'h000000003F07F87C00FE0001F801F02F03E000000063F618738E771BF1BF7C1C6FF8E0E1F0F07071FCE0381FDFB87E383871DE3B9DCEC7831FD871C638000000,
        char_line67 = 512'h000000001F01803F000000000003E03B07E000000077773C7B8E779BF1BF7F7E6FFCC3FBF1FDFCFDFDF87C1FDFB87EFEFEF3DE7B9DEECFC79FD9FDE6FE000000,
        char_line68 = 512'h000000000F81800FC0000000000FC00E07C00000003E773C7B8E77DBBBB07767630FC31B81DD8DCC73987C03183860CEC6FBDF7B9DEEDCC7871B9DF6E6000000,
        char_line69 = 512'h000000000FC00007F0000000003F00000F800000001C70366F8E77DBBB3F7F7E6387871DF1FF8EF871F07B831FB87EC1C7FBDFFB9DB6DC0DC71B8DF6FC000000,
        char_line70 = 512'h0000000007E00001FC00000000FE00001F000000001E707E6F8E77FB9F3F7F5F6387071FF1FB8E3C72F8FF031FB87CC7C7FEDFFB9DBEDCEFC71B8DFEBE000000,
        char_line71 = 512'h0000000003F000007F80000007F9E0003F0000000037707F678F777B9E3F7777638303BB81C1DDCC73B8EF031FBF7EEEEEEEDFFBBD9ECDDFC71BDDDEEE000000,
        char_line72 = 512'h0000000001F803381FF000007FE1E8007E0000000073F0E36787E73B8E3F777E638701F381C0F8FC71F07F831FBF7E7C7CEEDDB9F9DECFD8E719F9CE7C000000,
        char_line73 = 512'h0000000000FC037E07FFC01FFF83F800FC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line74 = 512'h00000000007E07FE00FFFFFFFC03F003F80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line75 = 512'h00000000003F87F8000FFFFFC003FC07F00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line76 = 512'h00000000001FC3FC0F003FF00303F00FC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line77 = 512'h00000000000FE0FC1F00000003E3783F800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line78 = 512'h000000000003F800FF07800601C0187F000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line79 = 512'h000000000001FE00FF0F9C3FC7F821FE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line80 = 512'h0000000000007F80FF8FF87FC7BC07F8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line81 = 512'h0000000000003FE0EC0FF07E01001FF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line82 = 512'h0000000000000FF8061FF07E07007FC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line83 = 512'h00000000000003FF000EF03E0603FF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line84 = 512'h00000000000000FFE000F01F001FFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line85 = 512'h000000000000003FFC00C00700FFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line86 = 512'h000000000000000FFFE000001FFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line87 = 512'h0000000000000001FFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line88 = 512'h00000000000000003FFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line89 = 512'h000000000000000003FFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line90 = 512'h0000000000000000001FFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line91 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line92 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line93 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line94 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line95 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line96 = 512'h0000000000000000000000000000000000000000000003F000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        char_line97 = 512'h00000000000000000000000000000000380000000000FFFE0000000001E00000000001C000000000000001800000000000000000000000000000000000000000,
        char_line98 = 512'h00000000000000000000000000000001FC000000000FFFFF8000000003F0070000000FF00000000000003FC000000000000F0000000000000000000000000000,
        char_line99 = 512'h0000000000000000000000000000003FFC000000003FF0FFE000000003F807C000003FF00000000000003FC000000000001F8000000000000000000000000000,
        char_line100 = 512'h000000000000000000000000000000FFF800000000FF800FF000000003FBC3E00001FFF000000000000007C000000000F80FC000000000000000000000000000,
        char_line101 = 512'h000000000000000000000000000000FFF00000000079C00FF800000001FFE1E0000FC3F00000000000000F8000000003FC0F8000000000000000000000000000,
        char_line102 = 512'h0000000000000000000000000000003FE00000000007E007F800000001FFF0E0000FE3C00000000000000F0000000003FC0F0000000000000000000000000000,
        char_line103 = 512'h0000000000000000000000000000008FDE000000F01FF007F800000001FFF0000007E7C00000000000000F7C00000001FE0F0000000000000000000000000000,
        char_line104 = 512'h00000000000000000000000000000387FE000001F03FF007F800000003FFF0000007F7800000000000001FFC00000001FE1F0000000000000000000000000000,
        char_line105 = 512'h000000000000000000000000000003CFFC000001F07FF007F000000003FFC0000007F7800000000000003FF800000000FE1E0000000000000000000000000000,
        char_line106 = 512'h000000000000000000000000000003EFF0000003F0FFF007F00000000FFF00000007F7800000000000003FF000000000FC7E0000000000000000000000000000,
        char_line107 = 512'h000000000000000000000000000007FFE3F00003F0FFE007F0000001FFF80000000FFFE0000000000000FF0000000000FFFF0000000000000000000000000000,
        char_line108 = 512'h000000000000000000000000000003FFFFF80003F0E7C003F0000003FFF00000000FFFF0000000000003FFC000000001FFFF0000000000000000000000000000,
        char_line109 = 512'h000000000000000000000000000001FFFFFC0007F00FF003F0000001FFF00000000FFFE000000000000FF9E00000001FFFFF0000000000000000000000000000,
        char_line110 = 512'h00000000000000000000000000000FFFFFFC0007F01FF003F0000000F9F3E000000FFFE000000000003FF0F80000001FFFFE0000000000000000000000000000,
        char_line111 = 512'h00000000000000000000000000003FFFE7F00007F07FF003F000000001F7E000000FFFC0000000000039F07C00001C0FFFFC0000000000000000000000000000,
        char_line112 = 512'h0000000000000000000000000000FFF19FE00007F0FFF003F000000001FFC000000FFFC0000000000001E03E00001E0FFFFE0000000000000000000000000000,
        char_line113 = 512'h0000000000000000000000000001FE03BF80000FF1FFF003E00000007FFF8000000FFFC0000000000003E03F80000E03F87F0000000000000000000000000000,
        char_line114 = 512'h0000000000000000000000000003E007FE00000FF1FFE003E0000001FFFF0000000FFFC0000000000003C01FC0000E03F3FE0000000000000000000000000000,
        char_line115 = 512'h0000000000000000000000000007C007F800000FF1FFC003E0000007FFFE00000007FFC0000000000007C06FFF800E03FFFC0000000000000000000000000000,
        char_line116 = 512'h000000000000000000000000000F800FF800000FF1FF9F03E000003FFFFC00000003FFFF80000000000FDFFFFFF80C01FFFC0000000000000000000000000000,
        char_line117 = 512'h000000000000000000000000001F803FE000000FF0FF1F03E000003FFFF80000000FFFFF80000000001FFFFFFFFC0007FC7C0000000000000000000000000000,
        char_line118 = 512'h000000000000000000000000001F00FF8000000FF0FF1F03E000003FFFF80000001EFFFF80000000007FFFCFFFFC003FF83C0000000000000000000000000000,
        char_line119 = 512'h000000000000000000000000001F01FEE000000FF1FFFE03E000001FFFF80000007FFFFE0000000000FFC700FFF800FFF03C0000000000000000000000000000,
        char_line120 = 512'h000000000000000000000000000C07FBF000000FF3FFFC03E0000001FFFE000000FFFFFC0000000001FE07F8780001F9F03C0000000000000000000000000000,
        char_line121 = 512'h00000000000000000000000000000FF3F000000FF7FFFC03E0000003E3FFC00003FFFFF00000000003FE0FF878000FC1E03C0000000000000000000000000000,
        char_line122 = 512'h00000000000000000000000000000FE0F000000FF7FFF803E0000007E1FFFC0003FFFFC07C0000007FFF3FF070000F81E03C0000000000000000000000000000,
        char_line123 = 512'h000000000000000000000000000003FEE000000FF7FFF003E000000FE1FFFFC003FFFFC0FC0000007FFF7FE0F0000FE0E03C0000000000000000000000000000,
        char_line124 = 512'h000000000000000000000000000007FFE000000FF3FE0003E000000FC1F87FFE00BFFFC0700000007FBF7F80E00003F0003C0000000000000000000000000000,
        char_line125 = 512'h00000000000000000000000000000FFFF000000FF1F00003F000001FFFF80FFFC07FFFC0000000007E3F0781E0000FF8007C0000000000000000000000000000,
        char_line126 = 512'h00000000000000000000000000000F1FFF00000FFFF80003F000003FFFF803FFC07FFFFC00000000183FF783C0007FFFFFF80000000000000000000000000000,
        char_line127 = 512'h00000000000000000000000000001E07FFE00007FFF00003F000007FFFF800FF8000FFFFE0000000003FFFC78001FFFFFFFFFFC0000000000000000000000000,
        char_line128 = 512'h00000000000000000000000000003C07FFFF0001FF800003F00000FE0FF8003F00000FFFFF800000001FFFE78001FFFFFFFFFFE0000000000000000000000000,
        char_line129 = 512'h00000000000000000000000000007007FFFFF8000000FE07F00000FC03F00000000000FFFFF80000001FFFFF0001FC3FFFFFFFE0000000000000000000000000,
        char_line130 = 512'h0000000000000000000000000000FFFC1FFFF8000000FFFFF00000F00000000000000007FFF80000001FFFFE00018000FFFFFFE0000000000000000000000000,
        char_line131 = 512'h0000000000000000000000000001FFF8073FF80000003FFFF000006000000000000000007FF80000001F87F80000000007FFFF00000000000000000000000000,
        char_line132 = 512'h000000000000000000000000000183F000000000000007FFC0000000000000000000000001F80000000000000000000000000000000000000000000000000000,
        char_line133 = 512'h00000000000000000000000000000000000000000000007F00000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // 图案显示逻辑
    wire display_active = (x_cnt >= 10'd180 && x_cnt < 10'd692) && (y_cnt >= 10'd190 && y_cnt <= 10'd323);
    reg [8:0] char_bit; // 用于行的每一列的位图

    // 在有效区域内显示图案
    always @(posedge clk_vga) begin
        if (!lcd_rst)
            char_bit <= 9'h1ff;
        else if (x_cnt == 10'd180)
            char_bit <= 9'd512;
        else if (display_active && x_cnt > 10'd180 && x_cnt < 10'd692)
            char_bit <= char_bit - 1'b1;
    end

    // 颜色输出逻辑
    reg [11:0] vga_rgb;
    always @ (posedge clk_vga) begin
        if (!lcd_rst || !display_active)
            vga_rgb <= 12'h000; // 黑色背景
        else begin
            case(y_cnt)
                10'd190:
                    if(char_line0[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd191:
                    if(char_line1[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd192:
                    if(char_line2[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd193:
                    if(char_line3[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd194:
                    if(char_line4[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd195:
                    if(char_line5[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd196:
                    if(char_line6[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd197:
                    if(char_line7[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd198:
                    if(char_line8[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd199:
                    if(char_line9[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd200:
                    if(char_line10[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd201:
                    if(char_line11[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd202:
                    if(char_line12[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd203:
                    if(char_line13[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd204:
                    if(char_line14[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd205:
                    if(char_line15[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd206:
                    if(char_line16[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd207:
                    if(char_line17[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd208:
                    if(char_line18[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd209:
                    if(char_line19[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd210:
                    if(char_line20[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd211:
                    if(char_line21[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd212:
                    if(char_line22[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd213:
                    if(char_line23[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd214:
                    if(char_line24[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd215:
                    if(char_line25[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd216:
                    if(char_line26[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd217:
                    if(char_line27[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd218:
                    if(char_line28[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd219:
                    if(char_line29[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd220:
                    if(char_line30[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd221:
                    if(char_line31[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd222:
                    if(char_line32[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd223:
                    if(char_line33[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd224:
                    if(char_line34[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd225:
                    if(char_line35[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd226:
                    if(char_line36[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd227:
                    if(char_line37[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd228:
                    if(char_line38[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd229:
                    if(char_line39[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd230:
                    if(char_line40[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd231:
                    if(char_line41[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd232:
                    if(char_line42[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd233:
                    if(char_line43[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd234:
                    if(char_line44[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd235:
                    if(char_line45[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd236:
                    if(char_line46[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd237:
                    if(char_line47[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd238:
                    if(char_line48[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd239:
                    if(char_line49[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd240:
                    if(char_line50[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd241:
                    if(char_line51[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd242:
                    if(char_line52[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd243:
                    if(char_line53[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd244:
                    if(char_line54[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd245:
                    if(char_line55[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd246:
                    if(char_line56[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd247:
                    if(char_line57[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd248:
                    if(char_line58[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd249:
                    if(char_line59[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd250:
                    if(char_line60[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd251:
                    if(char_line61[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd252:
                    if(char_line62[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd253:
                    if(char_line63[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd254:
                    if(char_line64[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd255:
                    if(char_line65[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd256:
                    if(char_line66[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd257:
                    if(char_line67[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd258:
                    if(char_line68[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd259:
                    if(char_line69[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd260:
                    if(char_line70[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd261:
                    if(char_line71[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd262:
                    if(char_line72[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd263:
                    if(char_line73[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd264:
                    if(char_line74[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd265:
                    if(char_line75[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd266:
                    if(char_line76[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd267:
                    if(char_line77[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd268:
                    if(char_line78[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd269:
                    if(char_line79[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd270:
                    if(char_line80[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd271:
                    if(char_line81[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd272:
                    if(char_line82[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd273:
                    if(char_line83[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd274:
                    if(char_line84[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd275:
                    if(char_line85[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd276:
                    if(char_line86[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd277:
                    if(char_line87[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd278:
                    if(char_line88[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd279:
                    if(char_line89[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd280:
                    if(char_line90[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd281:
                    if(char_line91[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd282:
                    if(char_line92[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd283:
                    if(char_line93[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd284:
                    if(char_line94[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd285:
                    if(char_line95[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd286:
                    if(char_line96[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd287:
                    if(char_line97[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd288:
                    if(char_line98[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd289:
                    if(char_line99[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd290:
                    if(char_line100[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd291:
                    if(char_line101[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd292:
                    if(char_line102[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd293:
                    if(char_line103[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd294:
                    if(char_line104[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd295:
                    if(char_line105[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd296:
                    if(char_line106[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd297:
                    if(char_line107[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd298:
                    if(char_line108[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd299:
                    if(char_line109[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd300:
                    if(char_line110[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd301:
                    if(char_line111[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd302:
                    if(char_line112[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd303:
                    if(char_line113[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd304:
                    if(char_line114[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd305:
                    if(char_line115[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd306:
                    if(char_line116[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd307:
                    if(char_line117[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd308:
                    if(char_line118[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd309:
                    if(char_line119[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd310:
                    if(char_line120[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd311:
                    if(char_line121[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd312:
                    if(char_line122[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd313:
                    if(char_line123[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd314:
                    if(char_line124[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd315:
                    if(char_line125[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd316:
                    if(char_line126[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd317:
                    if(char_line127[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd318:
                    if(char_line128[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd319:
                    if(char_line129[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd320:
                    if(char_line130[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd321:
                    if(char_line131[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd322:
                    if(char_line132[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd323:
                    if(char_line133[char_bit])
                        vga_rgb <=  12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                default:
                    vga_rgb <= 12'h000;
            endcase

        end
    end

    // 分配颜色输出
    assign vga_r = vga_rgb[11:8];
    assign vga_g = vga_rgb[7:4];
    assign vga_b = vga_rgb[3:0];

endmodule
