`define BLACK       12'b0000_0000_0000
module vga(
        input clk,               // 100MHz
        input lcd_rst,             // 复位信号
        input select,            // 模式选择
        output hsync,            // 行同步信号
        output vsync,            // 场同步信号
        output [3:0] vga_r,      // VGA红色信号
        output [3:0] vga_g,      // VGA绿色信号
        output [3:0] vga_b       // VGA蓝色信号
    );

    // 行和列计数
    reg [9:0] x_cnt;
    reg [9:0] y_cnt;
    reg clk_vga = 0;
    reg clk_cnt = 0;

    // 生成25MHz VGA时钟
    always @(posedge clk) begin
        if (!lcd_rst)
            clk_vga <= 0;
        else if (clk_cnt == 1) begin
            clk_vga <= ~clk_vga;
            clk_cnt <= 0;
        end
        else
            clk_cnt <= clk_cnt + 1;
    end

    // VGA行和列计数
    always @ (posedge clk_vga) begin
        if (!lcd_rst)
            x_cnt <= 10'd0;
        else if (x_cnt == 10'd799)
            x_cnt <= 10'd0;
        else
            x_cnt <= x_cnt + 1;
    end

    always @ (posedge clk_vga) begin
        if (!lcd_rst)
            y_cnt <= 10'd0;
        else if (x_cnt == 10'd799) begin
            if (y_cnt == 10'd524)
                y_cnt <= 10'd0;
            else
                y_cnt <= y_cnt + 1;
        end
    end

    // VGA同步信号生成
    reg hsync_r, vsync_r;
    always @ (posedge clk_vga) begin
        if (!lcd_rst)
            hsync_r <= 1'b1;
        else if (x_cnt == 10'd0)
            hsync_r <= 1'b0;
        else if (x_cnt == 10'd96)
            hsync_r <= 1'b1;
    end

    always @ (posedge clk_vga) begin
        if (!lcd_rst)
            vsync_r <= 1'b1;
        else if (y_cnt == 10'd0)
            vsync_r <= 1'b0;
        else if (y_cnt == 10'd2)
            vsync_r <= 1'b1;
    end

    assign hsync = hsync_r;
    assign vsync = vsync_r;

    // 定义图案数据
    //XUPT logo  512X256
    parameter

        char_line0 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line1 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line2 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line3 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line4 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line5 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line6 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line7 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line8 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line9 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line10 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line11 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line12 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line13 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line14 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line15 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line16 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line17 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line18 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line19 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line20 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line21 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line22 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line23 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line24 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line25 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line26 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line27 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line28 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line29 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line30 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line31 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line32 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line33 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line34 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line35 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line36 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line37 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line38 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line39 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line40 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line41 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line42 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line43 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line44 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line45 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line46 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line47 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line48 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line49 = 512'h0000000000000000000000000000000000000000000000000000000000001FFFFFE0000000000000000000000000000000000000000000000000000000000000,
    char_line50 = 512'h000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000,
    char_line51 = 512'h0000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000,
    char_line52 = 512'h00000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000,
    char_line53 = 512'h0000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000,
    char_line54 = 512'h00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000,
    char_line55 = 512'h0000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000,
    char_line56 = 512'h000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000,
    char_line57 = 512'h00000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000,
    char_line58 = 512'h0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000,
    char_line59 = 512'h000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000,
    char_line60 = 512'h00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000,
    char_line61 = 512'h0000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000,
    char_line62 = 512'h0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000,
    char_line63 = 512'h000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000,
    char_line64 = 512'h00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000,
    char_line65 = 512'h00000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000,
    char_line66 = 512'h0000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000,
    char_line67 = 512'h000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000,
    char_line68 = 512'h000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000,
    char_line69 = 512'h00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000,
    char_line70 = 512'h00000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000,
    char_line71 = 512'h0000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000,
    char_line72 = 512'h0000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000,
    char_line73 = 512'h000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000,
    char_line74 = 512'h000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000,
    char_line75 = 512'h00000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000,
    char_line76 = 512'h00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000,
    char_line77 = 512'h0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000,
    char_line78 = 512'h0000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000,
    char_line79 = 512'h0000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000,
    char_line80 = 512'h000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000,
    char_line81 = 512'h000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000,
    char_line82 = 512'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFF00000000000000000000000000000000,
    char_line83 = 512'h00000000000000000000000000000001FFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFF80000000000000000000000000000000,
    char_line84 = 512'h00000000000000000000000000000003FFFFFFFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000FFFFFFFFFFFC0000000000000000000000000000000,
    char_line85 = 512'h00000000000000000000000000000007FFFFFFFFFFE0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFFFFFFFE0000000000000000000000000000000,
    char_line86 = 512'h0000000000000000000000000000001FFFFFFFFFFFE00000003FFFFFFFFFFFFFFFFFFFFFFFFFFC00000007FFFFFFFFFFF8000000000000000000000000000000,
    char_line87 = 512'h0000000000000000000000000000003FFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFC000000000000000000000000000000,
    char_line88 = 512'h0000000000000000000000000000007FFFFFFFFFFFC0000000007FFFFFFFFC00003FFFFFFFFE0000000003FFFFFFFFFFFE000000000000000000000000000000,
    char_line89 = 512'h000000000000000000000000000000FFFFFFFFFFFF80000000000FFFFC0000000000003FFFF00000000001FFFFFFFFFFFF000000000000000000000000000000,
    char_line90 = 512'h000000000000000000000000000003FFFFFFFFFFFF800000000001F000000000000000000F800000000001FFFFFFFFFFFFC00000000000000000000000000000,
    char_line91 = 512'h000000000000000000000000000007FFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFE00000000000000000000000000000,
    char_line92 = 512'h000000000000000000000000000007FFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFE00000000000000000000000000000,
    char_line93 = 512'h00000000000000000000000000001FFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFF80000000000000000000000000000,
    char_line94 = 512'h00000000000000000000000000003FFFFFFFFFFFFF00000000000000000000000000000000000000000000FFFFFFFFFFFFFC0000000000000000000000000000,
    char_line95 = 512'h00000000000000000000000000003FFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFC0000000000000000000000000000,
    char_line96 = 512'h00000000000000000000000000007FFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFE0000000000000000000000000000,
    char_line97 = 512'h0000000000000000000000000000FFFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFF0000000000000000000000000000,
    char_line98 = 512'h0000000000000000000000000001FFFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFF8000000000000000000000000000,
    char_line99 = 512'h0000000000000000000000000003FFFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFFC000000000000000000000000000,
    char_line100 = 512'h0000000000000000000000000007FFFFFFFFFFFFFF80000000000000000000000000000000000000000003FFFFFFFFFFFFFFE000000000000000000000000000,
    char_line101 = 512'h000000000000000000000000000FFFFFFFFFFFFFFFC0000000000000000000000000000000000000000003FFFFFFFFFFFFFFF000000000000000000000000000,
    char_line102 = 512'h000000000000000000000000000FFFFFFFFFFFFFFFE0000000000000000000000000000000000000000007FFFFFFFFFFFFFFF000000000000000000000000000,
    char_line103 = 512'h000000000000000000000000001FFFFFFFFFFFFFFFE0000000000000000000000000000000000000000007FFFFFFFFFFFFFFF800000000000000000000000000,
    char_line104 = 512'h000000000000000000000000001FFFFFFFFFFFFFFFE0000000000000000000000000000000000000000007FFFFFFFFFFFFFFF800000000000000000000000000,
    char_line105 = 512'h000000000000000000000000003FFFFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFFFC00000000000000000000000000,
    char_line106 = 512'h000000000000000000000000007FFFFFFFFFFFFFFF00000000000000000000000000000000000000000000FFFFFFFFFFFFFFFE00000000000000000000000000,
    char_line107 = 512'h000000000000000000000000007FFFFFFFFFFFFFFC000000000000000000000000000000000000000000003FFFFFFFFFFFFFFE00000000000000000000000000,
    char_line108 = 512'h00000000000000000000000000FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000001FFFFFFFFFFFFFFF00000000000000000000000000,
    char_line109 = 512'h00000000000000000000000000FFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF00000000000000000000000000,
    char_line110 = 512'h00000000000000000000000001FFFFFFFFFFFFFFE00000000000000000000000000000000000000000000007FFFFFFFFFFFFFF80000000000000000000000000,
    char_line111 = 512'h00000000000000000000000003FFFFFFFFFFFFFFC00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFC0000000000000000000000000,
    char_line112 = 512'h00000000000000000000000003FFFFFFFFFFFFFF800000000000000000000000000000000000000000000001FFFFFFFFFFFFFFC0000000000000000000000000,
    char_line113 = 512'h00000000000000000000000003FFFFFFFFFFFFFF000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFC0000000000000000000000000,
    char_line114 = 512'h00000000000000000000000007FFFFFFFFFFFFFE0000000000000000000000000000000000000000000000007FFFFFFFFFFFFFE0000000000000000000000000,
    char_line115 = 512'h00000000000000000000000007FFFFFFFFFFFFFE0000000000000000000000000000000000000000000000007FFFFFFFFFFFFFE0000000000000000000000000,
    char_line116 = 512'h00000000000000000000000007FFFFFFFFFFFFFC0000000000000000000000000000000000000000000000003FFFFFFFFFFFFFE0000000000000000000000000,
    char_line117 = 512'h0000000000000000000000000FFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000003FFFFFFFFFFFFFF0000000000000000000000000,
    char_line118 = 512'h0000000000000000000000000FFFFFFFFFFFFFF80000000000000000000000000000000000000000000000001FFFFFFFFFFFFFF0000000000000000000000000,
    char_line119 = 512'h0000000000000000000000000FFFFFFFFFFFFFF80000000000000000000000000000000000000000000000001FFFFFFFFFFFFFF0000000000000000000000000,
    char_line120 = 512'h0000000000000000000000000FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFF0000000000000000000000000,
    char_line121 = 512'h0000000000000000000000001FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFF8000000000000000000000000,
    char_line122 = 512'h0000000000000000000000001FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFF8000000000000000000000000,
    char_line123 = 512'h0000000000000000000000001FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFF8000000000000000000000000,
    char_line124 = 512'h0000000000000000000000001FFFFFFFFFFFFFE000000000000000000000000000000000000000000000000007FFFFFFFFFFFFF8000000000000000000000000,
    char_line125 = 512'h0000000000000000000000001FFFFFFFFFFFFFE000000000000000000000000000000000000000000000000007FFFFFFFFFFFFF8000000000000000000000000,
    char_line126 = 512'h0000000000000000000000003FFFFFFFFFFFFFE000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFC000000000000000000000000,
    char_line127 = 512'h0000000000000000000000003FFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFF8000000000000000000000000,
    char_line128 = 512'h0000000000000000000000003FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFC000000000000000000000000,
    char_line129 = 512'h0000000000000000000000003FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFC000000000000000000000000,
    char_line130 = 512'h0000000000000000000000003FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFC000000000000000000000000,
    char_line131 = 512'h0000000000000000000000003FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFC000000000000000000000000,
    char_line132 = 512'h0000000000000000000000001FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFF8000000000000000000000000,
    char_line133 = 512'h0000000000000000000000003FFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFC000000000000000000000000,
    char_line134 = 512'h0000000000000000000000001FFFFFFFFFFFFFF80000000000000000000000000000000000000000000000001FFFFFFFFFFFFFF8000000000000000000000000,
    char_line135 = 512'h0000000000000000000000001FFFFFFFFFFFFFF80000000000000000000000000000000000000000000000001FFFFFFFFFFFFFF8000000000000000000000000,
    char_line136 = 512'h0000000000000000000000001FFFFFFFFFFFFFF80000000000000000000000000000000000000000000000001FFFFFFFFFFFFFF8000000000000000000000000,
    char_line137 = 512'h0000000000000000000000001FFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000003FFFFFFFFFFFFFF8000000000000000000000000,
    char_line138 = 512'h0000000000000000000000001FFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000003FFFFFFFFFFFFFF8000000000000000000000000,
    char_line139 = 512'h0000000000000000000000001FFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000007FFFFFFFFFFFFFF0000000000000000000000000,
    char_line140 = 512'h0000000000000000000000000FFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000007FFFFFFFFFFFFFF0000000000000000000000000,
    char_line141 = 512'h0000000000000000000000000FFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF0000000000000000000000000,
    char_line142 = 512'h0000000000000000000000000FFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFE0000000000000000000000000,
    char_line143 = 512'h00000000000000000000000007FFFFFFFFFFFFFF800000000000000000000000000000000000000000000001FFFFFFFFFFFFFFE0000000000000000000000000,
    char_line144 = 512'h00000000000000000000000007FFFFFFFFFFFFFFC00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFE0000000000000000000000000,
    char_line145 = 512'h00000000000000000000000007FFFFFFFFFFFFFFC00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFE0000000000000000000000000,
    char_line146 = 512'h00000000000000000000000003FFFFFFFFFFFFFFE00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFC0000000000000000000000000,
    char_line147 = 512'h00000000000000000000000003FFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFC0000000000000000000000000,
    char_line148 = 512'h00000000000000000000000001FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000001FFFFFFFFFFFFFFF80000000000000000000000000,
    char_line149 = 512'h00000000000000000000000001FFFFFFFFFFFFFFFC000000000000000000000000000000000000000000003FFFFFFFFFFFFFFF80000000000000000000000000,
    char_line150 = 512'h00000000000000000000000000FFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000FFFFFFFFFFFFFFFF00000000000000000000000000,
    char_line151 = 512'h00000000000000000000000000FFFFFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFFFF00000000000000000000000000,
    char_line152 = 512'h000000000000000000000000007FFFFFFFFFFFFFFFE0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFE00000000000000000000000000,
    char_line153 = 512'h000000000000000000000000007FFFFFFFFFFFFFFFF000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFE00000000000000000000000000,
    char_line154 = 512'h000000000000000000000000003FFFFFFFFFFFFFFFFC00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFC00000000000000000000000000,
    char_line155 = 512'h000000000000000000000000001FFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFF800000000000000000000000000,
    char_line156 = 512'h000000000000000000000000001FFFFFFFFFFFFFFFFFC000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF800000000000000000000000000,
    char_line157 = 512'h000000000000000000000000000FFFFFFFFFFFFFFFFFF80000000000000000000000000000000000001FFFFFFFFFFFFFFFFFF000000000000000000000000000,
    char_line158 = 512'h000000000000000000000000000FFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFE000000000000000000000000000,
    char_line159 = 512'h0000000000000000000000000007FFFFFFFFFFFFFFFFFFE00000000000000000000000000000000007FFFFFFFFFFFFFFFFFFE000000000000000000000000000,
    char_line160 = 512'h0000000000000000000000000003FFFFFFFFFFFFFFFFFFFC000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFC000000000000000000000000000,
    char_line161 = 512'h0000000000000000000000000001FFFFFFFF83FFFFFFFFFFC0000000000000000000000000000007FFFFFFFFFFFFFFFFFFFF8000000000000000000000000000,
    char_line162 = 512'h0000000000000000000000000000FFFFFFF0000FFFFFFFFFFE00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000,
    char_line163 = 512'h00000000000000000000000000007FFFFFF80001FFFFFFFFFFF80000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000,
    char_line164 = 512'h00000000000000000000000000003FFFFFFC00003FFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000,
    char_line165 = 512'h00000000000000000000000000001FFFFFFF000007FFFFFFFFFFFFFF8000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000,
    char_line166 = 512'h00000000000000000000000000001FFFFFFFE00001FFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000,
    char_line167 = 512'h00000000000000000000000000000FFFFFFFFC0000FFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000,
    char_line168 = 512'h000000000000000000000000000003FFFFFFFF00003FFFFFFFFFFFFE00000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000,
    char_line169 = 512'h000000000000000000000000000001FFFFFFFFC0001FFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000,
    char_line170 = 512'h000000000000000000000000000000FFFFFFFFE0000FFFFFFFFFFFF800000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000,
    char_line171 = 512'h0000000000000000000000000000007FFFFFFFF80003FFFFFFFFFFF000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000,
    char_line172 = 512'h0000000000000000000000000000003FFFFFFFFC0001FFFFFFFFFFE0000000000000000007FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000,
    char_line173 = 512'h0000000000000000000000000000001FFFFFFFFE00007FFFFFFFFFE0000000000000000007FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000,
    char_line174 = 512'h00000000000000000000000000000007FFFFFFFF00001FFFFFFFFFC0000000000000000003FFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000,
    char_line175 = 512'h00000000000000000000000000000003FFFFFFFF800007FFFFFFFFC0000000000000000003FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000,
    char_line176 = 512'h00000000000000000000000000000001FFFFFFFFC00000FFFFFFFF80000000000000000001FFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000,
    char_line177 = 512'h000000000000000000000000000000007FFFFFFFE000000FFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000,
    char_line178 = 512'h000000000000000000000000000000003FFFFFFFF00000000FC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000,
    char_line179 = 512'h000000000000000000000000000000001FFFFFFFF800000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000,
    char_line180 = 512'h0000000000000000000000000000000007FFFFFFFC00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000,
    char_line181 = 512'h0000000000000000000000000000000001FFFFFFFE00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000,
    char_line182 = 512'h0000000000000000000000000000000000FFFFFFFF00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000,
    char_line183 = 512'h00000000000000000000000000000000003FFFFFFFC0000000000000000000000000000001FFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000,
    char_line184 = 512'h00000000000000000000000000000000000FFFFFFFF0000000000000000000000000000001FFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000,
    char_line185 = 512'h000000000000000000000000000000000007FFFFFFFC000000000000000000000000000001FFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000,
    char_line186 = 512'h000000000000000000000000000000000001FFFFFFFF800000000000000000000000000001FFFFFFFFFFFFFFFFFF000000000000000000000000000000000000,
    char_line187 = 512'h0000000000000000000000000000000000007FFFFFFFF00000000000000000000000000001FFFFFFFFFFFFFFFFFE000000000000000000000000000000000000,
    char_line188 = 512'h0000000000000000000000000000000000001FFFFFFFFF8000000000000000000000000001FFFFFFFFFFFFFFFFF0000000000000000000000000000000000000,
    char_line189 = 512'h00000000000000000000000000000000000007FFFFFFFFFE00001F80000000000000000001FFFFFFFFFFFFFFFFE0000000000000000000000000000000000000,
    char_line190 = 512'h00000000000000000000000000000000000000FFFFFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFFFF00000000000000000000000000000000000000,
    char_line191 = 512'h000000000000000000000000000000000000003FFFFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFFFC00000000000000000000000000000000000000,
    char_line192 = 512'h000000000000000000000000000000000000000FFFFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFFF000000000000000000000000000000000000000,
    char_line193 = 512'h0000000000000000000000000000000000000003FFFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFF8000000000000000000000000000000000000000,
    char_line194 = 512'h00000000000000000000000000000000000000007FFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFE0000000000000000000000000000000000000000,
    char_line195 = 512'h00000000000000000000000000000000000000000FFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFF00000000000000000000000000000000000000000,
    char_line196 = 512'h000000000000000000000000000000000000000003FFFFFFFFFFFF80000000000000000001FFFFFFFFFFFF800000000000000000000000000000000000000000,
    char_line197 = 512'h0000000000000000000000000000000000000000003FFFFFFFFFFF80000000000000000001FFFFFFFFFFFC000000000000000000000000000000000000000000,
    char_line198 = 512'h00000000000000000000000000000000000000000007FFFFFFFFFF80000000000000000001FFFFFFFFFFF0000000000000000000000000000000000000000000,
    char_line199 = 512'h00000000000000000000000000000000000000000000FFFFFFFFFF80000000000000000001FFFFFFFFFF00000000000000000000000000000000000000000000,
    char_line200 = 512'h000000000000000000000000000000000000000000001FFFFFFFFF80000000000000000001FFFFFFFFF800000000000000000000000000000000000000000000,
    char_line201 = 512'h0000000000000000000000000000000000000000000001FFFFFFFF80000000000000000001FFFFFFFF8000000000000000000000000000000000000000000000,
    char_line202 = 512'h00000000000000000000000000000000000000000000001FFFFFFF80000000000000000001FFFFFFF80000000000000000000000000000000000000000000000,
    char_line203 = 512'h000000000000000000000000000000000000000000000001FFFFFF80000000000000000001FFFFFF800000000000000000000000000000000000000000000000,
    char_line204 = 512'h0000000000000000000000000000000000000000000000001FFFFF00000000000000000000FFFFF8000000000000000000000000000000000000000000000000,
    char_line205 = 512'h00000000000000000000000000000000000000000000000000FFFE000000000000000000007FFF00000000000000000000000000000000000000000000000000,
    char_line206 = 512'h0000000000000000000000000000000000000000000000000003F0000000000000000000000FE000000000000000000000000000000000000000000000000000,
    char_line207 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line208 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line209 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line210 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line211 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line212 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line213 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line214 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line215 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line216 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line217 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line218 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line219 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line220 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line221 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line222 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line223 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line224 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line225 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line226 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line227 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line228 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line229 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line230 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line231 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line232 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line233 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line234 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line235 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line236 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line237 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line238 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line239 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line240 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line241 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line242 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line243 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line244 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line245 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line246 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line247 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line248 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line249 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line250 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line251 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line252 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line253 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line254 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    char_line255 = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // 图案显示逻辑
    wire display_active = (x_cnt >= 10'd180 && x_cnt < 10'd692) && (y_cnt >= 10'd190 && y_cnt <= 10'd445);
    reg [8:0] char_bit; // 用于行的每一列的位图

    // 在有效区域内显示图案
    always @(posedge clk_vga) begin
        if (!lcd_rst)
            char_bit <= 9'h1ff;
        else if (x_cnt == 10'd180)
            char_bit <= 9'd512;
        else if (display_active && x_cnt > 10'd180 && x_cnt < 10'd692)
            char_bit <= char_bit - 1'b1;
    end

    // 颜色输出逻辑
    reg [11:0] vga_rgb;
    always @ (posedge clk_vga) begin
        if (!lcd_rst || !display_active)
            vga_rgb <= 12'h000; // 黑色背景
        else begin
            case(y_cnt)
                10'd190:
                    if(char_line0[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd191:
                    if(char_line1[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd192:
                    if(char_line2[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd193:
                    if(char_line3[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd194:
                    if(char_line4[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd195:
                    if(char_line5[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd196:
                    if(char_line6[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd197:
                    if(char_line7[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd198:
                    if(char_line8[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd199:
                    if(char_line9[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd200:
                    if(char_line10[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd201:
                    if(char_line11[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd202:
                    if(char_line12[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd203:
                    if(char_line13[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd204:
                    if(char_line14[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd205:
                    if(char_line15[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd206:
                    if(char_line16[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd207:
                    if(char_line17[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd208:
                    if(char_line18[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd209:
                    if(char_line19[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd210:
                    if(char_line20[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd211:
                    if(char_line21[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd212:
                    if(char_line22[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd213:
                    if(char_line23[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd214:
                    if(char_line24[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd215:
                    if(char_line25[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd216:
                    if(char_line26[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd217:
                    if(char_line27[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd218:
                    if(char_line28[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd219:
                    if(char_line29[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd220:
                    if(char_line30[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd221:
                    if(char_line31[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd222:
                    if(char_line32[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd223:
                    if(char_line33[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd224:
                    if(char_line34[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd225:
                    if(char_line35[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd226:
                    if(char_line36[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd227:
                    if(char_line37[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd228:
                    if(char_line38[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd229:
                    if(char_line39[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd230:
                    if(char_line40[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd231:
                    if(char_line41[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd232:
                    if(char_line42[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd233:
                    if(char_line43[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd234:
                    if(char_line44[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd235:
                    if(char_line45[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd236:
                    if(char_line46[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd237:
                    if(char_line47[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd238:
                    if(char_line48[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd239:
                    if(char_line49[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd240:
                    if(char_line50[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd241:
                    if(char_line51[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd242:
                    if(char_line52[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd243:
                    if(char_line53[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd244:
                    if(char_line54[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd245:
                    if(char_line55[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd246:
                    if(char_line56[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd247:
                    if(char_line57[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd248:
                    if(char_line58[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd249:
                    if(char_line59[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd250:
                    if(char_line60[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd251:
                    if(char_line61[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd252:
                    if(char_line62[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd253:
                    if(char_line63[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd254:
                    if(char_line64[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd255:
                    if(char_line65[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd256:
                    if(char_line66[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd257:
                    if(char_line67[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd258:
                    if(char_line68[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd259:
                    if(char_line69[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd260:
                    if(char_line70[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd261:
                    if(char_line71[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd262:
                    if(char_line72[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd263:
                    if(char_line73[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd264:
                    if(char_line74[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd265:
                    if(char_line75[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd266:
                    if(char_line76[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd267:
                    if(char_line77[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd268:
                    if(char_line78[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd269:
                    if(char_line79[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd270:
                    if(char_line80[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd271:
                    if(char_line81[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd272:
                    if(char_line82[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd273:
                    if(char_line83[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd274:
                    if(char_line84[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd275:
                    if(char_line85[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd276:
                    if(char_line86[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd277:
                    if(char_line87[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd278:
                    if(char_line88[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd279:
                    if(char_line89[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd280:
                    if(char_line90[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd281:
                    if(char_line91[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd282:
                    if(char_line92[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd283:
                    if(char_line93[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd284:
                    if(char_line94[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd285:
                    if(char_line95[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd286:
                    if(char_line96[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd287:
                    if(char_line97[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd288:
                    if(char_line98[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd289:
                    if(char_line99[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd290:
                    if(char_line100[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd291:
                    if(char_line101[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd292:
                    if(char_line102[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd293:
                    if(char_line103[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd294:
                    if(char_line104[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd295:
                    if(char_line105[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd296:
                    if(char_line106[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd297:
                    if(char_line107[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd298:
                    if(char_line108[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd299:
                    if(char_line109[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd300:
                    if(char_line110[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd301:
                    if(char_line111[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd302:
                    if(char_line112[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd303:
                    if(char_line113[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd304:
                    if(char_line114[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd305:
                    if(char_line115[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd306:
                    if(char_line116[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd307:
                    if(char_line117[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd308:
                    if(char_line118[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd309:
                    if(char_line119[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd310:
                    if(char_line120[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd311:
                    if(char_line121[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd312:
                    if(char_line122[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd313:
                    if(char_line123[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd314:
                    if(char_line124[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd315:
                    if(char_line125[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd316:
                    if(char_line126[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd317:
                    if(char_line127[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd318:
                    if(char_line128[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd319:
                    if(char_line129[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd320:
                    if(char_line130[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd321:
                    if(char_line131[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd322:
                    if(char_line132[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd323:
                    if(char_line133[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd324:
                    if(char_line134[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd325:
                    if(char_line135[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd326:
                    if(char_line136[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd327:
                    if(char_line137[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd328:
                    if(char_line138[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd329:
                    if(char_line139[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd330:
                    if(char_line140[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd331:
                    if(char_line141[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd332:
                    if(char_line142[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd333:
                    if(char_line143[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd334:
                    if(char_line144[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd335:
                    if(char_line145[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd336:
                    if(char_line146[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd337:
                    if(char_line147[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd338:
                    if(char_line148[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd339:
                    if(char_line149[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd340:
                    if(char_line150[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd341:
                    if(char_line151[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd342:
                    if(char_line152[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd343:
                    if(char_line153[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd344:
                    if(char_line154[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd345:
                    if(char_line155[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd346:
                    if(char_line156[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd347:
                    if(char_line157[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd348:
                    if(char_line158[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd349:
                    if(char_line159[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd350:
                    if(char_line160[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd351:
                    if(char_line161[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd352:
                    if(char_line162[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd353:
                    if(char_line163[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd354:
                    if(char_line164[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd355:
                    if(char_line165[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd356:
                    if(char_line166[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd357:
                    if(char_line167[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd358:
                    if(char_line168[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd359:
                    if(char_line169[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd360:
                    if(char_line170[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd361:
                    if(char_line171[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd362:
                    if(char_line172[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd363:
                    if(char_line173[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd364:
                    if(char_line174[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd365:
                    if(char_line175[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd366:
                    if(char_line176[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd367:
                    if(char_line177[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd368:
                    if(char_line178[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd369:
                    if(char_line179[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd370:
                    if(char_line180[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd371:
                    if(char_line181[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd372:
                    if(char_line182[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd373:
                    if(char_line183[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd374:
                    if(char_line184[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd375:
                    if(char_line185[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd376:
                    if(char_line186[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd377:
                    if(char_line187[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd378:
                    if(char_line188[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd379:
                    if(char_line189[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd380:
                    if(char_line190[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd381:
                    if(char_line191[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd382:
                    if(char_line192[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd383:
                    if(char_line193[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd384:
                    if(char_line194[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd385:
                    if(char_line195[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd386:
                    if(char_line196[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd387:
                    if(char_line197[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd388:
                    if(char_line198[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd389:
                    if(char_line199[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd390:
                    if(char_line200[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd391:
                    if(char_line201[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd392:
                    if(char_line202[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd393:
                    if(char_line203[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd394:
                    if(char_line204[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd395:
                    if(char_line205[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd396:
                    if(char_line206[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd397:
                    if(char_line207[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd398:
                    if(char_line208[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd399:
                    if(char_line209[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd400:
                    if(char_line210[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd401:
                    if(char_line211[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd402:
                    if(char_line212[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd403:
                    if(char_line213[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd404:
                    if(char_line214[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd405:
                    if(char_line215[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd406:
                    if(char_line216[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd407:
                    if(char_line217[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd408:
                    if(char_line218[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd409:
                    if(char_line219[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd410:
                    if(char_line220[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd411:
                    if(char_line221[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd412:
                    if(char_line222[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd413:
                    if(char_line223[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd414:
                    if(char_line224[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd415:
                    if(char_line225[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd416:
                    if(char_line226[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd417:
                    if(char_line227[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd418:
                    if(char_line228[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd419:
                    if(char_line229[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd420:
                    if(char_line230[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd421:
                    if(char_line231[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd422:
                    if(char_line232[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd423:
                    if(char_line233[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd424:
                    if(char_line234[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd425:
                    if(char_line235[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd426:
                    if(char_line236[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd427:
                    if(char_line237[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd428:
                    if(char_line238[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd429:
                    if(char_line239[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd430:
                    if(char_line240[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd431:
                    if(char_line241[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd432:
                    if(char_line242[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd433:
                    if(char_line243[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd434:
                    if(char_line244[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd435:
                    if(char_line245[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd436:
                    if(char_line246[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd437:
                    if(char_line247[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd438:
                    if(char_line248[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd439:
                    if(char_line249[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd440:
                    if(char_line250[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd441:
                    if(char_line251[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd442:
                    if(char_line252[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd443:
                    if(char_line253[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd444:
                    if(char_line254[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                10'd445:
                    if(char_line255[char_bit])
                        vga_rgb <= 12'd1111_1111_1111;
                    else
                        vga_rgb <= `BLACK;
                default:
                    vga_rgb <= 12'h000;
            endcase

        end
    end

    // 分配颜色输出
    assign vga_r = vga_rgb[11:8];
    assign vga_g = vga_rgb[7:4];
    assign vga_b = vga_rgb[3:0];

endmodule
